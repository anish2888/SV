//dff
